// test bench for input activation controller

`timescale 1ns/1ps
module tb_weight_in_ctrl();


endmodule
