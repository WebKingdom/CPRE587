// test bench for input activation controller

`timescale 1ns/1ps
module tb_input_act_ctrl();


endmodule
